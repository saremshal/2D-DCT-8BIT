`timescale 1ns / 1ps


module tbStimVerify(

    );
endmodule
